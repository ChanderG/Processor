//Data Memory

//???


module dataMemory();








endmodule
