//Meta level

//One level above the Processor

//Will create processor and feed clock from here

module topLevel();

